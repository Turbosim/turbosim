// this module includes compilaiton flags wich controls simulation or compilation
`ifndef _compilation_flags
`define _compilation_flags

// switch this flags on / off according to working mode (simmulation / synthesis)
//`define SYNTHESIS
`define SIMULATION


`endif