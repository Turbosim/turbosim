// DATA derived from module add1 !!!!!!!!!!!!!!!!
// table may be used turbo sim to hold the cell functionality delay and connectivity
// table width is 88 bits
// where first 4 bits holds the primitive type
// next is 16 bits that holds the primitive delay in ps
// next is 12 bits the holds the net index of the output pin - pin0 bit 11 is set if exist
// next is 16 bits for 4 input nets:
// 	12 bits the holds the net index of the input pin  - pinX bit 11 is set if exist
// 	4 bits that holds the input pin current value, set to x, R/W field
0_0327_871_84e_2_000_3_000_3_000_3    //    0 U10     |  not    807 ps   n24    n140    x UC      z UC      z UC      z 
5_019e_833_811_2_834_2_000_3_000_3    //    1 U100    |  nand   414 ps   n116   b[10]   x n117    x UC      z UC      z 
5_030c_834_835_2_836_2_000_3_000_3    //    2 U101    |  nand   780 ps   n117   n118    x n119    x UC      z UC      z 
2_0510_84e_84f_2_850_2_000_3_000_3    //    3 U102    |  and   1296 ps   n140   n141    x n142    x UC      z UC      z 
5_069c_84f_80b_2_879_2_000_3_000_3    //    4 U103    |  nand  1692 ps   n141   a[5]    x n31     x UC      z UC      z 
5_0511_850_81b_2_851_2_000_3_000_3    //    5 U104    |  nand  1297 ps   n142   b[5]    x n143    x UC      z UC      z 
5_04d1_851_852_2_87d_2_000_3_000_3    //    6 U105    |  nand  1233 ps   n143   n144    x n35     x UC      z UC      z 
2_0314_8c0_826_2_827_2_000_3_000_3    //    7 U106    |  and    788 ps   n96    n104    x n105    x UC      z UC      z 
5_00bb_826_802_2_82b_2_000_3_000_3    //    8 U107    |  nand   187 ps   n104   a[11]   x n109    x UC      z UC      z 
5_015a_827_812_2_828_2_000_3_000_3    //    9 U108    |  nand   346 ps   n105   b[11]   x n106    x UC      z UC      z 
5_00a2_828_829_2_82a_2_000_3_000_3    //   10 U109    |  nand   162 ps   n106   n107    x n108    x UC      z UC      z 
0_00b3_869_849_2_000_3_000_3_000_3    //   11 U11     |  not    179 ps   n17    n136    x UC      z UC      z UC      z 
2_02eb_849_84a_2_84b_2_000_3_000_3    //   12 U110    |  and    747 ps   n136   n137    x n138    x UC      z UC      z 
5_0484_84a_80c_2_871_2_000_3_000_3    //   13 U111    |  nand  1156 ps   n137   a[6]    x n24     x UC      z UC      z 
5_0675_84b_81c_2_84c_2_000_3_000_3    //   14 U112    |  nand  1653 ps   n138   b[6]    x n139    x UC      z UC      z 
5_053a_84c_84e_2_875_2_000_3_000_3    //   15 U113    |  nand  1338 ps   n139   n140    x n28     x UC      z UC      z 
2_02cc_8b4_8bd_2_8be_2_000_3_000_3    //   16 U114    |  and    716 ps   n85    n93     x n94     x UC      z UC      z 
5_0194_8bd_803_2_8c2_2_000_3_000_3    //   17 U115    |  nand   404 ps   n93    a[12]   x n98     x UC      z UC      z 
5_05e8_8be_813_2_8bf_2_000_3_000_3    //   18 U116    |  nand  1512 ps   n94    b[12]   x n95     x UC      z UC      z 
5_06d8_8bf_8c0_2_8c1_2_000_3_000_3    //   19 U117    |  nand  1752 ps   n95    n96     x n97     x UC      z UC      z 
2_0444_845_846_2_847_2_000_3_000_3    //   20 U118    |  and   1092 ps   n132   n133    x n134    x UC      z UC      z 
5_0655_846_80d_2_869_2_000_3_000_3    //   21 U119    |  nand  1621 ps   n133   a[7]    x n17     x UC      z UC      z 
0_0756_821_845_2_000_3_000_3_000_3    //   22 U12     |  not   1878 ps   n10    n132    x UC      z UC      z UC      z 
5_04b1_847_81d_2_848_2_000_3_000_3    //   23 U120    |  nand  1201 ps   n134   b[7]    x n135    x UC      z UC      z 
5_05f9_848_849_2_86e_2_000_3_000_3    //   24 U121    |  nand  1529 ps   n135   n136    x n21     x UC      z UC      z 
2_0286_8a5_8b1_2_8b2_2_000_3_000_3    //   25 U122    |  and    646 ps   n71    n82     x n83     x UC      z UC      z 
5_0056_8b1_804_2_8b6_2_000_3_000_3    //   26 U123    |  nand    86 ps   n82    a[13]   x n87     x UC      z UC      z 
5_0462_8b2_814_2_8b3_2_000_3_000_3    //   27 U124    |  nand  1122 ps   n83    b[13]   x n84     x UC      z UC      z 
5_06ce_8b3_8b4_2_8b5_2_000_3_000_3    //   28 U125    |  nand  1742 ps   n84    n85     x n86     x UC      z UC      z 
2_012e_835_83e_2_83f_2_000_3_000_3    //   29 U126    |  and    302 ps   n118   n126    x n127    x UC      z UC      z 
5_0619_83f_81f_2_840_2_000_3_000_3    //   30 U127    |  nand  1561 ps   n127   b[9]    x n128    x UC      z UC      z 
5_055a_83e_80f_2_877_2_000_3_000_3    //   31 U128    |  nand  1370 ps   n126   a[9]    x n3      x UC      z UC      z 
3_03c5_840_877_2_80f_2_000_3_000_3    //   32 U129    |  or     965 ps   n128   n3      x a[9]    x UC      z UC      z 
0_0050_82b_829_2_000_3_000_3_000_3    //   33 U13     |  not     80 ps   n109   n107    x UC      z UC      z UC      z 
5_02fa_8a0_8a8_2_8a9_2_000_3_000_3    //   34 U130    |  nand   762 ps   n67    n74     x n75     x UC      z UC      z 
3_0697_8a8_8aa_2_816_2_000_3_000_3    //   35 U131    |  or    1687 ps   n74    n76     x b[15]   x UC      z UC      z 
5_0319_8a9_816_2_8aa_2_000_3_000_3    //   36 U132    |  nand   793 ps   n75    b[15]   x n76     x UC      z UC      z 
0_015c_8aa_806_2_000_3_000_3_000_3    //   37 U133    |  not    348 ps   n76    a[15]   x UC      z UC      z UC      z 
5_0200_893_818_2_894_2_000_3_000_3    //   38 U134    |  nand   512 ps   n55    b[2]    x n56     x UC      z UC      z 
5_00c8_88b_819_2_88c_2_000_3_000_3    //   39 U135    |  nand   200 ps   n48    b[3]    x n49     x UC      z UC      z 
5_063a_884_81a_2_885_2_000_3_000_3    //   40 U136    |  nand  1594 ps   n41    b[4]    x n42     x UC      z UC      z 
5_002a_87c_81b_2_87d_2_000_3_000_3    //   41 U137    |  nand    42 ps   n34    b[5]    x n35     x UC      z UC      z 
5_0703_874_81c_2_875_2_000_3_000_3    //   42 U138    |  nand  1795 ps   n27    b[6]    x n28     x UC      z UC      z 
5_04f7_86d_81d_2_86e_2_000_3_000_3    //   43 U139    |  nand  1271 ps   n20    b[7]    x n21     x UC      z UC      z 
0_016a_8c2_8c0_2_000_3_000_3_000_3    //   44 U14     |  not    362 ps   n98    n96     x UC      z UC      z UC      z 
5_0616_842_81e_2_84d_2_000_3_000_3    //   45 U140    |  nand  1558 ps   n13    b[8]    x n14     x UC      z UC      z 
5_0317_83d_811_2_836_2_000_3_000_3    //   46 U141    |  nand   791 ps   n125   b[10]   x n119    x UC      z UC      z 
5_0449_831_812_2_82a_2_000_3_000_3    //   47 U142    |  nand  1097 ps   n114   b[11]   x n108    x UC      z UC      z 
5_0128_825_813_2_8c1_2_000_3_000_3    //   48 U143    |  nand   296 ps   n103   b[12]   x n97     x UC      z UC      z 
5_03b0_8bc_814_2_8b5_2_000_3_000_3    //   49 U144    |  nand   944 ps   n92    b[13]   x n86     x UC      z UC      z 
5_05d2_8b0_815_2_8a6_2_000_3_000_3    //   50 U145    |  nand  1490 ps   n81    b[14]   x n72     x UC      z UC      z 
5_06b7_89b_817_2_89c_2_000_3_000_3    //   51 U146    |  nand  1719 ps   n62    b[1]    x n63     x UC      z UC      z 
5_01ac_8a2_815_2_8a4_2_000_3_000_3    //   52 U147    |  nand   428 ps   n69    b[14]   x n70     x UC      z UC      z 
5_007b_8a4_8a5_2_8a6_2_000_3_000_3    //   53 U148    |  nand   123 ps   n70    n71     x n72     x UC      z UC      z 
5_020d_8a1_805_2_8a7_2_000_3_000_3    //   54 U149    |  nand   525 ps   n68    a[14]   x n73     x UC      z UC      z 
0_05ca_8b6_8b4_2_000_3_000_3_000_3    //   55 U15     |  not   1482 ps   n87    n85     x UC      z UC      z UC      z 
0_03de_894_808_2_000_3_000_3_000_3    //   56 U150    |  not    990 ps   n56    a[2]    x UC      z UC      z UC      z 
0_04a3_88c_809_2_000_3_000_3_000_3    //   57 U151    |  not   1187 ps   n49    a[3]    x UC      z UC      z UC      z 
0_03f4_885_80a_2_000_3_000_3_000_3    //   58 U152    |  not   1012 ps   n42    a[4]    x UC      z UC      z UC      z 
0_06be_87d_80b_2_000_3_000_3_000_3    //   59 U153    |  not   1726 ps   n35    a[5]    x UC      z UC      z UC      z 
0_069c_875_80c_2_000_3_000_3_000_3    //   60 U154    |  not   1692 ps   n28    a[6]    x UC      z UC      z UC      z 
0_01b6_86e_80d_2_000_3_000_3_000_3    //   61 U155    |  not    438 ps   n21    a[7]    x UC      z UC      z UC      z 
0_0177_84d_80e_2_000_3_000_3_000_3    //   62 U156    |  not    375 ps   n14    a[8]    x UC      z UC      z UC      z 
0_02c5_836_801_2_000_3_000_3_000_3    //   63 U157    |  not    709 ps   n119   a[10]   x UC      z UC      z UC      z 
0_00fa_82a_802_2_000_3_000_3_000_3    //   64 U158    |  not    250 ps   n108   a[11]   x UC      z UC      z UC      z 
0_004a_8c1_803_2_000_3_000_3_000_3    //   65 U159    |  not     74 ps   n97    a[12]   x UC      z UC      z UC      z 
0_0524_8a7_8a5_2_000_3_000_3_000_3    //   66 U16     |  not   1316 ps   n73    n71     x UC      z UC      z UC      z 
0_002d_8b5_804_2_000_3_000_3_000_3    //   67 U160    |  not     45 ps   n86    a[13]   x UC      z UC      z UC      z 
0_01cb_8a6_805_2_000_3_000_3_000_3    //   68 U161    |  not    459 ps   n72    a[14]   x UC      z UC      z UC      z 
5_04e7_898_81f_2_8a3_2_000_3_000_3    //   69 U162    |  nand  1255 ps   n6     b[9]    x n7      x UC      z UC      z 
0_02ad_89c_807_2_000_3_000_3_000_3    //   70 U163    |  not    685 ps   n63    a[1]    x UC      z UC      z UC      z 
0_008c_865_810_2_000_3_000_3_000_3    //   71 U164    |  not    140 ps   n161   b[0]    x UC      z UC      z UC      z 
0_0790_866_800_2_000_3_000_3_000_3    //   72 U165    |  not   1936 ps   n162   a[0]    x UC      z UC      z UC      z 
5_0376_8c4_867_2_868_2_000_3_000_3    //   73 U166    |  nand   886 ps   o[0]   n163    x n164    x UC      z UC      z 
5_061c_867_800_2_865_2_000_3_000_3    //   74 U167    |  nand  1564 ps   n163   a[0]    x n161    x UC      z UC      z 
5_0145_868_810_2_866_2_000_3_000_3    //   75 U168    |  nand   325 ps   n164   b[0]    x n162    x UC      z UC      z 
3_0219_89a_89c_2_817_2_000_3_000_3    //   76 U169    |  or     537 ps   n61    n63     x b[1]    x UC      z UC      z 
0_07a4_838_835_2_000_3_000_3_000_3    //   77 U17     |  not   1956 ps   n120   n118    x UC      z UC      z UC      z 
3_030b_892_894_2_818_2_000_3_000_3    //   78 U170    |  or     779 ps   n54    n56     x b[2]    x UC      z UC      z 
3_0529_88a_88c_2_819_2_000_3_000_3    //   79 U171    |  or    1321 ps   n47    n49     x b[3]    x UC      z UC      z 
3_04a6_883_885_2_81a_2_000_3_000_3    //   80 U172    |  or    1190 ps   n40    n42     x b[4]    x UC      z UC      z 
3_00d2_87b_87d_2_81b_2_000_3_000_3    //   81 U173    |  or     210 ps   n33    n35     x b[5]    x UC      z UC      z 
3_039e_873_875_2_81c_2_000_3_000_3    //   82 U174    |  or     926 ps   n26    n28     x b[6]    x UC      z UC      z 
3_05b0_86b_86e_2_81d_2_000_3_000_3    //   83 U175    |  or    1456 ps   n19    n21     x b[7]    x UC      z UC      z 
3_0323_837_84d_2_81e_2_000_3_000_3    //   84 U176    |  or     803 ps   n12    n14     x b[8]    x UC      z UC      z 
3_0033_88d_8a3_2_81f_2_000_3_000_3    //   85 U177    |  or      51 ps   n5     n7      x b[9]    x UC      z UC      z 
3_0481_83c_836_2_811_2_000_3_000_3    //   86 U178    |  or    1153 ps   n124   n119    x b[10]   x UC      z UC      z 
3_00b1_830_82a_2_812_2_000_3_000_3    //   87 U179    |  or     177 ps   n113   n108    x b[11]   x UC      z UC      z 
4_05a9_8cc_88e_2_88f_2_000_3_000_3    //   88 U18     |  nor   1449 ps   o[2]   n50     x n51     x UC      z UC      z 
3_01f5_824_8c1_2_813_2_000_3_000_3    //   89 U180    |  or     501 ps   n102   n97     x b[12]   x UC      z UC      z 
3_0494_8bb_8b5_2_814_2_000_3_000_3    //   90 U181    |  or    1172 ps   n91    n86     x b[13]   x UC      z UC      z 
3_06c9_8af_8a6_2_815_2_000_3_000_3    //   91 U182    |  or    1737 ps   n80    n72     x b[14]   x UC      z UC      z 
0_0310_8a3_80f_2_000_3_000_3_000_3    //   92 U183    |  not    784 ps   n7     a[9]    x UC      z UC      z UC      z 
2_00e1_88f_890_2_891_2_000_3_000_3    //   93 U19     |  and    225 ps   n51    n52     x n53     x UC      z UC      z 
4_0286_88e_890_2_891_2_000_3_000_3    //   94 U20     |  nor    646 ps   n50    n52     x n53     x UC      z UC      z 
5_0250_891_892_2_893_2_000_3_000_3    //   95 U21     |  nand   592 ps   n53    n54     x n55     x UC      z UC      z 
4_06e2_8cd_886_2_887_2_000_3_000_3    //   96 U22     |  nor   1762 ps   o[3]   n43     x n44     x UC      z UC      z 
2_014b_887_888_2_889_2_000_3_000_3    //   97 U23     |  and    331 ps   n44    n45     x n46     x UC      z UC      z 
4_0044_886_888_2_889_2_000_3_000_3    //   98 U24     |  nor     68 ps   n43    n45     x n46     x UC      z UC      z 
5_01d2_889_88a_2_88b_2_000_3_000_3    //   99 U25     |  nand   466 ps   n46    n47     x n48     x UC      z UC      z 
4_065c_8ce_87e_2_87f_2_000_3_000_3    //  100 U26     |  nor   1628 ps   o[4]   n36     x n37     x UC      z UC      z 
2_0217_87f_880_2_881_2_000_3_000_3    //  101 U27     |  and    535 ps   n37    n38     x n39     x UC      z UC      z 
4_04dc_87e_880_2_881_2_000_3_000_3    //  102 U28     |  nor   1244 ps   n36    n38     x n39     x UC      z UC      z 
5_07ce_881_883_2_884_2_000_3_000_3    //  103 U29     |  nand  1998 ps   n39    n40     x n41     x UC      z UC      z 
4_023a_8cf_876_2_878_2_000_3_000_3    //  104 U30     |  nor    570 ps   o[5]   n29     x n30     x UC      z UC      z 
2_03a1_878_879_2_87a_2_000_3_000_3    //  105 U31     |  and    929 ps   n30    n31     x n32     x UC      z UC      z 
4_0386_876_879_2_87a_2_000_3_000_3    //  106 U32     |  nor    902 ps   n29    n31     x n32     x UC      z UC      z 
5_03e2_87a_87b_2_87c_2_000_3_000_3    //  107 U33     |  nand   994 ps   n32    n33     x n34     x UC      z UC      z 
4_00d2_8d0_86f_2_870_2_000_3_000_3    //  108 U34     |  nor    210 ps   o[6]   n22     x n23     x UC      z UC      z 
2_0208_870_871_2_872_2_000_3_000_3    //  109 U35     |  and    520 ps   n23    n24     x n25     x UC      z UC      z 
4_0589_86f_871_2_872_2_000_3_000_3    //  110 U36     |  nor   1417 ps   n22    n24     x n25     x UC      z UC      z 
5_0472_872_873_2_874_2_000_3_000_3    //  111 U37     |  nand  1138 ps   n25    n26     x n27     x UC      z UC      z 
4_0039_8d1_858_2_863_2_000_3_000_3    //  112 U38     |  nor     57 ps   o[7]   n15     x n16     x UC      z UC      z 
2_0061_863_869_2_86a_2_000_3_000_3    //  113 U39     |  and     97 ps   n16    n17     x n18     x UC      z UC      z 
0_03f2_899_864_2_000_3_000_3_000_3    //  114 U4      |  not   1010 ps   n60    n160    x UC      z UC      z UC      z 
4_05b1_858_869_2_86a_2_000_3_000_3    //  115 U40     |  nor   1457 ps   n15    n17     x n18     x UC      z UC      z 
5_0141_86a_86b_2_86d_2_000_3_000_3    //  116 U41     |  nand   321 ps   n18    n19     x n20     x UC      z UC      z 
4_06e3_8d2_8ae_2_8b9_2_000_3_000_3    //  117 U42     |  nor   1763 ps   o[8]   n8      x n9      x UC      z UC      z 
2_06c5_8b9_821_2_82c_2_000_3_000_3    //  118 U43     |  and   1733 ps   n9     n10     x n11     x UC      z UC      z 
4_02d9_8ae_821_2_82c_2_000_3_000_3    //  119 U44     |  nor    729 ps   n8     n10     x n11     x UC      z UC      z 
5_027d_82c_837_2_842_2_000_3_000_3    //  120 U45     |  nand   637 ps   n11    n12     x n13     x UC      z UC      z 
4_0184_8d3_820_2_86c_2_000_3_000_3    //  121 U46     |  nor    388 ps   o[9]   n1      x n2      x UC      z UC      z 
2_04c8_86c_877_2_882_2_000_3_000_3    //  122 U47     |  and   1224 ps   n2     n3      x n4      x UC      z UC      z 
4_077a_820_877_2_882_2_000_3_000_3    //  123 U48     |  nor   1914 ps   n1     n3      x n4      x UC      z UC      z 
5_034f_882_88d_2_898_2_000_3_000_3    //  124 U49     |  nand   847 ps   n4     n5      x n6      x UC      z UC      z 
4_0598_864_865_2_866_2_000_3_000_3    //  125 U5      |  nor   1432 ps   n160   n161    x n162    x UC      z UC      z 
4_00fd_8c5_839_2_83a_2_000_3_000_3    //  126 U50     |  nor    253 ps   o[10]  n121    x n122    x UC      z UC      z 
2_0311_83a_838_2_83b_2_000_3_000_3    //  127 U51     |  and    785 ps   n122   n120    x n123    x UC      z UC      z 
4_0721_839_838_2_83b_2_000_3_000_3    //  128 U52     |  nor   1825 ps   n121   n120    x n123    x UC      z UC      z 
5_046c_83b_83c_2_83d_2_000_3_000_3    //  129 U53     |  nand  1132 ps   n123   n124    x n125    x UC      z UC      z 
4_0794_8c6_82d_2_82e_2_000_3_000_3    //  130 U54     |  nor   1940 ps   o[11]  n110    x n111    x UC      z UC      z 
2_0135_82e_82b_2_82f_2_000_3_000_3    //  131 U55     |  and    309 ps   n111   n109    x n112    x UC      z UC      z 
4_0372_82d_82b_2_82f_2_000_3_000_3    //  132 U56     |  nor    882 ps   n110   n109    x n112    x UC      z UC      z 
5_03ac_82f_830_2_831_2_000_3_000_3    //  133 U57     |  nand   940 ps   n112   n113    x n114    x UC      z UC      z 
4_07c5_8c7_8c3_2_822_2_000_3_000_3    //  134 U58     |  nor   1989 ps   o[12]  n99     x n100    x UC      z UC      z 
2_01fc_822_8c2_2_823_2_000_3_000_3    //  135 U59     |  and    508 ps   n100   n98     x n101    x UC      z UC      z 
0_0784_890_85f_2_000_3_000_3_000_3    //  136 U6      |  not   1924 ps   n52    n156    x UC      z UC      z UC      z 
4_03a8_8c3_8c2_2_823_2_000_3_000_3    //  137 U60     |  nor    936 ps   n99    n98     x n101    x UC      z UC      z 
5_06d4_823_824_2_825_2_000_3_000_3    //  138 U61     |  nand  1748 ps   n101   n102    x n103    x UC      z UC      z 
4_0755_8c8_8b7_2_8b8_2_000_3_000_3    //  139 U62     |  nor   1877 ps   o[13]  n88     x n89     x UC      z UC      z 
2_00f5_8b8_8b6_2_8ba_2_000_3_000_3    //  140 U63     |  and    245 ps   n89    n87     x n90     x UC      z UC      z 
4_0212_8b7_8b6_2_8ba_2_000_3_000_3    //  141 U64     |  nor    530 ps   n88    n87     x n90     x UC      z UC      z 
5_0604_8ba_8bb_2_8bc_2_000_3_000_3    //  142 U65     |  nand  1540 ps   n90    n91     x n92     x UC      z UC      z 
4_071a_8c9_8ab_2_8ac_2_000_3_000_3    //  143 U66     |  nor   1818 ps   o[14]  n77     x n78     x UC      z UC      z 
2_0559_8ac_8a7_2_8ad_2_000_3_000_3    //  144 U67     |  and   1369 ps   n78    n73     x n79     x UC      z UC      z 
4_0667_8ab_8a7_2_8ad_2_000_3_000_3    //  145 U68     |  nor   1639 ps   n77    n73     x n79     x UC      z UC      z 
5_033a_8ad_8af_2_8b0_2_000_3_000_3    //  146 U69     |  nand   826 ps   n79    n80     x n81     x UC      z UC      z 
0_0154_888_85b_2_000_3_000_3_000_3    //  147 U7      |  not    340 ps   n45    n152    x UC      z UC      z UC      z 
4_07ad_8ca_89d_2_89e_2_000_3_000_3    //  148 U70     |  nor   1965 ps   o[15]  n64     x n65     x UC      z UC      z 
2_0553_89e_89f_2_8a0_2_000_3_000_3    //  149 U71     |  and   1363 ps   n65    n66     x n67     x UC      z UC      z 
4_03c9_89d_8a0_2_89f_2_000_3_000_3    //  150 U72     |  nor    969 ps   n64    n67     x n66     x UC      z UC      z 
5_03ef_89f_8a1_2_8a2_2_000_3_000_3    //  151 U73     |  nand  1007 ps   n66    n68     x n69     x UC      z UC      z 
5_0239_8cb_895_2_896_2_000_3_000_3    //  152 U74     |  nand   569 ps   o[1]   n57     x n58     x UC      z UC      z 
3_046c_896_897_2_899_2_000_3_000_3    //  153 U75     |  or    1132 ps   n58    n59     x n60     x UC      z UC      z 
5_0747_895_897_2_899_2_000_3_000_3    //  154 U76     |  nand  1863 ps   n57    n59     x n60     x UC      z UC      z 
5_0382_897_89a_2_89b_2_000_3_000_3    //  155 U77     |  nand   898 ps   n59    n61     x n62     x UC      z UC      z 
5_0671_877_841_2_843_2_000_3_000_3    //  156 U78     |  nand  1649 ps   n3     n129    x n130    x UC      z UC      z 
5_00da_841_80e_2_821_2_000_3_000_3    //  157 U79     |  nand   218 ps   n129   a[8]    x n10     x UC      z UC      z 
0_0398_880_856_2_000_3_000_3_000_3    //  158 U8      |  not    920 ps   n38    n148    x UC      z UC      z UC      z 
5_075f_843_81e_2_844_2_000_3_000_3    //  159 U80     |  nand  1887 ps   n130   b[8]    x n131    x UC      z UC      z 
5_00e2_844_845_2_84d_2_000_3_000_3    //  160 U81     |  nand   226 ps   n131   n132    x n14     x UC      z UC      z 
2_06da_85f_860_2_861_2_000_3_000_3    //  161 U82     |  and   1754 ps   n156   n157    x n158    x UC      z UC      z 
5_030a_861_817_2_862_2_000_3_000_3    //  162 U83     |  nand   778 ps   n158   b[1]    x n159    x UC      z UC      z 
5_0095_860_807_2_864_2_000_3_000_3    //  163 U84     |  nand   149 ps   n157   a[1]    x n160    x UC      z UC      z 
5_077a_862_89c_2_899_2_000_3_000_3    //  164 U85     |  nand  1914 ps   n159   n63     x n60     x UC      z UC      z 
2_016d_85b_85c_2_85d_2_000_3_000_3    //  165 U86     |  and    365 ps   n152   n153    x n154    x UC      z UC      z 
5_0273_85c_808_2_890_2_000_3_000_3    //  166 U87     |  nand   627 ps   n153   a[2]    x n52     x UC      z UC      z 
5_0593_85d_818_2_85e_2_000_3_000_3    //  167 U88     |  nand  1427 ps   n154   b[2]    x n155    x UC      z UC      z 
5_07a5_85e_85f_2_894_2_000_3_000_3    //  168 U89     |  nand  1957 ps   n155   n156    x n56     x UC      z UC      z 
0_00c5_879_852_2_000_3_000_3_000_3    //  169 U9      |  not    197 ps   n31    n144    x UC      z UC      z UC      z 
2_05e1_856_857_2_859_2_000_3_000_3    //  170 U90     |  and   1505 ps   n148   n149    x n150    x UC      z UC      z 
5_0295_857_809_2_888_2_000_3_000_3    //  171 U91     |  nand   661 ps   n149   a[3]    x n45     x UC      z UC      z 
5_0482_859_819_2_85a_2_000_3_000_3    //  172 U92     |  nand  1154 ps   n150   b[3]    x n151    x UC      z UC      z 
5_02cf_85a_85b_2_88c_2_000_3_000_3    //  173 U93     |  nand   719 ps   n151   n152    x n49     x UC      z UC      z 
2_045e_852_853_2_854_2_000_3_000_3    //  174 U94     |  and   1118 ps   n144   n145    x n146    x UC      z UC      z 
5_03c4_853_80a_2_880_2_000_3_000_3    //  175 U95     |  nand   964 ps   n145   a[4]    x n38     x UC      z UC      z 
5_0148_854_81a_2_855_2_000_3_000_3    //  176 U96     |  nand   328 ps   n146   b[4]    x n147    x UC      z UC      z 
5_01b6_855_856_2_885_2_000_3_000_3    //  177 U97     |  nand   438 ps   n147   n148    x n42     x UC      z UC      z 
2_06f1_829_832_2_833_2_000_3_000_3    //  178 U98     |  and   1777 ps   n107   n115    x n116    x UC      z UC      z 
5_03a2_832_801_2_838_2_000_3_000_3    //  179 U99     |  nand   930 ps   n115   a[10]   x n120    x UC      z UC      z 
