`timescale 1ns /1ps

module add4 ( o, a, b );
  output [15:0] o;
  input [15:0] a;
  input [15:0] b;
  wire   n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163,
         n164;
	
  wire   a0,a1, a2, a3, a4, a5, a6, a7,
         a8, a9, a10, a11, a12, a13,
         a14, a15;
		 
  wire   b0,b1, b2, b3, b4, b5, b6, b7,
         b8, b9, b10, b11, b12, b13,
         b14, b15;
		 
  wire   o0,o1, o2, o3, o4, o5, o6, o7,
         o8, o9, o10, o11, o12, o13,
         o14, o15;
		 
		 
  buf	#(0.716) G0 ( a0, a[0]);
  buf	#(0.716) G1 ( a1, a[0]);
  buf	#(0.716) G2 ( a2, a[1]); 
  buf	#(0.716) G3 ( a3, a[1]);
  buf	#(0.716) G4 ( a4, a[2]);
  buf	#(0.716) G5 ( a5, a[2]);
  buf	#(0.716) G6 ( a6, a[3]); 
  buf	#(0.716) G7 ( a7, a[3]);
  buf	#(0.716) G8 ( a8, a[4]);
  buf	#(0.716) G9 ( a9, a[4]);
  buf	#(0.716) G10 ( a10, a[5]); 
  buf	#(0.716) G11 ( a11, a[5]);
  buf	#(0.716) G12 ( a12, a[6]);
  buf	#(0.716) G13 ( a13, a[6]);
  buf	#(0.716) G14 ( a14, a[7]); 
  buf	#(0.716) G15 ( a15, a[7]);
  
   buf	#(0.716) H0 ( b0, b[0]);
  buf	#(0.716) H1 ( b1, b[0]);
  buf	#(0.716) H2 ( b2, b[1]); 
  buf	#(0.716) H3 ( b3, b[1]);
  buf	#(0.716) H4 ( b4, b[2]);
  buf	#(0.716) H5 ( b5, b[2]);
  buf	#(0.716) H6 ( b6, b[3]); 
  buf	#(0.716) H7 ( b7, b[3]);
  buf	#(0.716) H8 ( b8, b[4]);
  buf	#(0.716) H9 ( b9, b[4]);
  buf	#(0.716) H10 ( b10, b[5]); 
  buf	#(0.716) H11 ( b11, b[5]);
  buf	#(0.716) H12 ( b12, b[6]);
  buf	#(0.716) H13 ( b13, b[6]);
  buf	#(0.716) H14 ( b14, b[7]); 
  buf	#(0.716) H15 ( b15, b[7]);
                           
  nand  #(0.716) K0  ( o[0],o0,o1,o2,o3);
  nand  #(0.716) K1  ( o[1],o4,o5,o6,o7);
  nand  #(0.716) K2  ( o[2],o8,o9,o10,o11);
  nand  #(0.716) K3  ( o[3],o12,o13,o14,o15);
  
                     
  
  
  
  


  not	#(1.000) U4 ( n60, n160 );
  nor	#(1.000) U5 ( n160, n161, n162 );
  not	#(1.000) U6 ( n52, n156 );
  not	#(1.000) U7 ( n45, n152 );
  not	#(1.000) U8 ( n38, n148 );
  not	#(1.000) U9 ( n31, n144 );
  not	#(1.000) U10 ( n24, n140 );
  not	#(1.000) U11 ( n17, n136 );
  not	#(1.000) U12 ( n10, n132 );
  not	#(1.000) U13 ( n109, n107 );
  not	#(1.000) U14 ( n98, n96 );
  not	#(1.000) U15 ( n87, n85 );
  not	#(1.000) U16 ( n73, n71 );
  not	#(1.000) U17 ( n120, n118 );
  nor	#(1.000) U18 ( o2, n50, n51 );
  and	#(1.000) U19 ( n51, n52, n53 );
  nor	#(1.000) U20 ( n50, n52, n53 );
  nand	#(1.000) U21 ( n53, n54, n55 );
  nor	#(1.000) U22 ( o3, n43, n44 );
  and	#(1.000) U23 ( n44, n45, n46 );
  nor	#(1.000) U24 ( n43, n45, n46 );
  nand	#(1.000) U25 ( n46, n47, n48 );
  nor	#(1.000) U26 ( o4, n36, n37 );
  and	#(1.000) U27 ( n37, n38, n39 );
  nor	#(1.000) U28 ( n36, n38, n39 );
  nand	#(1.000) U29 ( n39, n40, n41 );
  nor	#(1.000) U30 ( o5, n29, n30 );
  and	#(1.000) U31 ( n30, n31, n32 );
  nor	#(1.000) U32 ( n29, n31, n32 );
  nand	#(1.000) U33 ( n32, n33, n34 );
  nor	#(1.000) U34 ( o6, n22, n23 );
  and	#(1.000) U35 ( n23, n24, n25 );
  nor	#(1.000) U36 ( n22, n24, n25 );
  nand	#(1.000) U37 ( n25, n26, n27 );
  nor	#(1.000) U38 ( o7, n15, n16 );
  and	#(1.000) U39 ( n16, n17, n18 );
  nor	#(1.000) U40 ( n15, n17, n18 );
  nand	#(1.000) U41 ( n18, n19, n20 );
  nor	#(1.000) U42 ( o8, n8, n9 );
  and	#(1.000) U43 ( n9, n10, n11 );
  nor	#(1.000) U44 ( n8, n10, n11 );
  nand	#(1.000) U45 ( n11, n12, n13 );
  nor	#(1.000) U46 ( o9, n1, n2 );
  and	#(1.000) U47 ( n2, n3, n4 );
  nor	#(1.000) U48 ( n1, n3, n4 );
  nand	#(1.000) U49 ( n4, n5, n6 );
  nor	#(1.000) U50 ( o10, n121, n122 );
  and	#(1.000) U51 ( n122, n120, n123 );
  nor	#(1.000) U52 ( n121, n120, n123 );
  nand	#(1.000) U53 ( n123, n124, n125 );
  nor	#(1.000) U54 ( o11, n110, n111 );
  and	#(1.000) U55 ( n111, n109, n112 );
  nor	#(1.000) U56 ( n110, n109, n112 );
  nand	#(1.000) U57 ( n112, n113, n114 );
  nor	#(1.000) U58 ( o12, n99, n100 );
  and	#(1.000) U59 ( n100, n98, n101 );
  nor	#(1.000) U60 ( n99, n98, n101 );
  nand	#(1.000) U61 ( n101, n102, n103 );
  nor	#(1.000) U62 ( o13, n88, n89 );
  and	#(1.000) U63 ( n89, n87, n90 );
  nor	#(1.000) U64 ( n88, n87, n90 );
  nand	#(1.000) U65 ( n90, n91, n92 );
  nor	#(1.000) U66 ( o14, n77, n78 );
  and	#(1.000) U67 ( n78, n73, n79 );
  nor	#(1.000) U68 ( n77, n73, n79 );
  nand	#(1.000) U69 ( n79, n80, n81 );
  nor	#(1.000) U70 ( o15, n64, n65 );
  and	#(1.000) U71 ( n65, n66, n67 );
  nor	#(1.000) U72 ( n64, n67, n66 );
  nand	#(1.000) U73 ( n66, n68, n69 );
  nand	#(1.000) U74 ( o1, n57, n58 );
  or	#(1.000) U75 ( n58, n59, n60 );
  nand	#(1.000) U76 ( n57, n59, n60 );
  nand	#(1.000) U77 ( n59, n61, n62 );
  nand	#(1.000) U78 ( n3, n129, n130 );
  nand	#(1.000) U79 ( n129, a8, n10 );
  nand	#(1.000) U80 ( n130, b8, n131 );
  nand	#(1.000) U81 ( n131, n132, n14 );
  and	#(1.000) U82 ( n156, n157, n158 );
  nand	#(1.000) U83 ( n158, b1, n159 );
  nand	#(1.000) U84 ( n157, a1, n160 );
  nand	#(1.000) U85 ( n159, n63, n60 );
  and	#(1.000) U86 ( n152, n153, n154 );
  nand	#(1.000) U87 ( n153, a2, n52 );
  nand	#(1.000) U88 ( n154, b2, n155 );
  nand	#(1.000) U89 ( n155, n156, n56 );
  and	#(1.000) U90 ( n148, n149, n150 );
  nand	#(1.000) U91 ( n149, a3, n45 );
  nand	#(1.000) U92 ( n150, b3, n151 );
  nand	#(1.000) U93 ( n151, n152, n49 );
  and	#(1.000) U94 ( n144, n145, n146 );
  nand	#(1.000) U95 ( n145, a4, n38 );
  nand	#(1.000) U96 ( n146, b4, n147 );
  nand	#(1.000) U97 ( n147, n148, n42 );
  and	#(1.000) U98 ( n107, n115, n116 );
  nand	#(1.000) U99 ( n115, a10, n120 );
  nand	#(1.000) U100 ( n116, b10, n117 );
  nand	#(1.000) U101 ( n117, n118, n119 );
  and	#(1.000) U102 ( n140, n141, n142 );
  nand	#(1.000) U103 ( n141, a5, n31 );
  nand	#(1.000) U104 ( n142, b5, n143 );
  nand	#(1.000) U105 ( n143, n144, n35 );
  and	#(1.000) U106 ( n96, n104, n105 );
  nand	#(1.000) U107 ( n104, a11, n109 );
  nand	#(1.000) U108 ( n105, b11, n106 );
  nand	#(1.000) U109 ( n106, n107, n108 );
  and	#(1.000) U110 ( n136, n137, n138 );
  nand	#(1.000) U111 ( n137, a6, n24 );
  nand	#(1.000) U112 ( n138, b6, n139 );
  nand	#(1.000) U113 ( n139, n140, n28 );
  and	#(1.000) U114 ( n85, n93, n94 );
  nand	#(1.000) U115 ( n93, a12, n98 );
  nand	#(1.000) U116 ( n94, b12, n95 );
  nand	#(1.000) U117 ( n95, n96, n97 );
  and	#(1.000) U118 ( n132, n133, n134 );
  nand	#(1.000) U119 ( n133, a7, n17 );
  nand	#(1.000) U120 ( n134, b7, n135 );
  nand	#(1.000) U121 ( n135, n136, n21 );
  and	#(1.000) U122 ( n71, n82, n83 );
  nand	#(1.000) U123 ( n82, a13, n87 );
  nand	#(1.000) U124 ( n83, b13, n84 );
  nand	#(1.000) U125 ( n84, n85, n86 );
  and	#(1.000) U126 ( n118, n126, n127 );
  nand	#(1.000) U127 ( n127, b9, n128 );
  nand	#(1.000) U128 ( n126, a9, n3 );
  or	#(1.000) U129 ( n128, n3, a9 );
  nand	#(1.000) U130 ( n67, n74, n75 );
  or	#(1.000) U131 ( n74, n76, b15 );
  nand	#(1.000) U132 ( n75, b15, n76 );
  not	#(1.000) U133 ( n76, a15 );
  nand	#(1.000) U134 ( n55, b2, n56 );
  nand	#(1.000) U135 ( n48, b3, n49 );
  nand	#(1.000) U136 ( n41, b4, n42 );
  nand	#(1.000) U137 ( n34, b5, n35 );
  nand	#(1.000) U138 ( n27, b6, n28 );
  nand	#(1.000) U139 ( n20, b7, n21 );
  nand	#(1.000) U140 ( n13, b8, n14 );
  nand	#(1.000) U141 ( n125, b10, n119 );
  nand	#(1.000) U142 ( n114, b11, n108 );
  nand	#(1.000) U143 ( n103, b12, n97 );
  nand	#(1.000) U144 ( n92, b13, n86 );
  nand	#(1.000) U145 ( n81, b14, n72 );
  nand	#(1.000) U146 ( n62, b1, n63 );
  nand	#(1.000) U147 ( n69, b14, n70 );
  nand	#(1.000) U148 ( n70, n71, n72 );
  nand	#(1.000) U149 ( n68, a14, n73 );
  not	#(1.000) U150 ( n56, a2 );
  not	#(1.000) U151 ( n49, a3 );
  not	#(1.000) U152 ( n42, a4 );
  not	#(1.000) U153 ( n35, a5 );
  not	#(1.000) U154 ( n28, a6 );
  not	#(1.000) U155 ( n21, a7 );
  not	#(1.000) U156 ( n14, a8 );
  not	#(1.000) U157 ( n119, a10 );
  not	#(1.000) U158 ( n108, a11 );
  not	#(1.000) U159 ( n97, a12 );
  not	#(1.000) U160 ( n86, a13 );
  not	#(1.000) U161 ( n72, a14 );
  nand	#(1.000) U162 ( n6, b9, n7 );
  not	#(1.000) U163 ( n63, a1 );
  not	#(1.000) U164 ( n161, b0 );
  not	#(1.000) U165 ( n162, a0 );
  nand	#(1.000) U166 ( o0, n163, n164 );
  nand	#(1.000) U167 ( n163, a0, n161 );
  nand	#(1.000) U168 ( n164, b0, n162 );
  or	#(1.000) U169 ( n61, n63, b1 );
  or	#(1.000) U170 ( n54, n56, b2 );
  or	#(1.000) U171 ( n47, n49, b3 );
  or	#(1.000) U172 ( n40, n42, b4 );
  or	#(1.000) U173 ( n33, n35, b5 );
  or	#(1.000) U174 ( n26, n28, b6 );
  or	#(1.000) U175 ( n19, n21, b7 );
  or	#(1.000) U176 ( n12, n14, b8 );
  or	#(1.000) U177 ( n5, n7, b9 );
  or	#(1.000) U178 ( n124, n119, b10 );
  or	#(1.000) U179 ( n113, n108, b11 );
  or	#(1.000) U180 ( n102, n97, b12 );
  or	#(1.000) U181 ( n91, n86, b13 );
  or	#(1.000) U182 ( n80, n72, b14 );
  not	#(1.000) U183 ( n7, a9 );
  
  wire   d1, d2, d3, d4, d5, d6, d7,
         d8, d9, d10, d11, d12, d13,
         d14, d15, d16, d17, d18, d19,
         d20, d21, d22, d23, d24, d25,
         d26, d27, d28, d29, d30, d31,
         d32, d33, d34, d35, d36, d37,
         d38, d39, d40, d41, d42, d43,
         d44, d45, d46, d47, d48, d49,
         d50, d51, d52, d53, d54, d55,
         d56, d57, d58, d59, d60, d61,
         d62, d63, d64, d65, d66, d67,
         d68, d69, d70, d71, d72, d73,
         d74, d75, d76, d77, d78, d79,
         d80, d81, d82, d83, d84, d85,
         d86, d87, d88, d89, d90, d91,
         d92, d93, d94, d95, d96, d97,
         d98, d99, d100, d101, d102, d103,
         d104, d105, d106, d107, d108,
         d109, d110, d111, d112, d113,
         d114, d115, d116, d117, d118,
         d119, d120, d121, d122, d123,
         d124, d125, d126, d127, d128,
         d129, d130, d131, d132, d133,
         d134, d135, d136, d137, d138,
         d139, d140, d141, d142, d143,
         d144, d145, d146, d147, d148,
         d149, d150, d151, d152, d153,
         d154, d155, d156, d157, d158,
         d159, d160, d161, d162, d163,
         d164;
	
  wire   c0,c1, c2, c3, c4, c5, c6, c7,
         c8, c9, c10, c11, c12, c13,
         c14, c15;
		 
  wire   e0,e1, e2, e3, e4, e5, e6, e7,
         e8, e9, e10, e11, e12, e13,
         e14, e15;
		 
  wire   f0,f1, f2, f3, f4, f5, f6, f7,
         f8, f9, f10, f11, f12, f13,
         f14, f15;
		 
		 
  buf	#(0.716) GW0 ( c0, a[0]);
  buf	#(0.716) GW1 ( c1, a[0]);
  buf	#(0.716) GW2 ( c2, a[1]); 
  buf	#(0.716) GW3 ( c3, a[1]);
  buf	#(0.716) GW4 ( c4, a[2]);
  buf	#(0.716) GW5 ( c5, a[2]);
  buf	#(0.716) GW6 ( c6, a[3]); 
  buf	#(0.716) GW7 ( c7, a[3]);
  buf	#(0.716) GW8 ( c8, a[4]);
  buf	#(0.716) GW9 ( c9, a[4]);
  buf	#(0.716) GW10 ( c10, a[5]); 
  buf	#(0.716) GW11 ( c11, a[5]);
  buf	#(0.716) GW12 ( c12, a[6]);
  buf	#(0.716) GW13 ( c13, a[6]);
  buf	#(0.716) GW14 ( c14, a[7]); 
  buf	#(0.716) GW15 ( c15, a[7]);
  
   buf	#(0.716) HW0 ( e0, b[0]);
  buf	#(0.716) HW1 ( e1, b[0]);
  buf	#(0.716) HW2 ( e2, b[1]); 
  buf	#(0.716) HW3 ( e3, b[1]);
  buf	#(0.716) HW4 ( e4, b[2]);
  buf	#(0.716) HW5 ( e5, b[2]);
  buf	#(0.716) HW6 ( e6, b[3]); 
  buf	#(0.716) HW7 ( e7, b[3]);
  buf	#(0.716) HW8 ( e8, b[4]);
  buf	#(0.716) HW9 ( e9, b[4]);
  buf	#(0.716) HW10 ( e10, b[5]); 
  buf	#(0.716) HW11 ( e11, b[5]);
  buf	#(0.716) HW12 ( e12, b[6]);
  buf	#(0.716) HW13 ( e13, b[6]);
  buf	#(0.716) HW14 ( e14, b[7]); 
  buf	#(0.716) HW15 ( e15, b[7]);
                               
  nand  #(0.716) KW0  ( o[4],f0,f1,f2,f3);
  nand  #(0.716) KW1  ( o[5],f4,f5,f6,f7);
  nand  #(0.716) KW2  ( o[6],f8,f9,f10,f11);
  nand  #(0.716) KW3  ( o[7],f12,f13,f14,f15);
  
                     
  
  
  
  


  not	#(1.000) UW4 ( d60, d160 );
  nor	#(1.000) UW5 ( d160, d161, d162 );
  not	#(1.000) UW6 ( d52, d156 );
  not	#(1.000) UW7 ( d45, d152 );
  not	#(1.000) UW8 ( d38, d148 );
  not	#(1.000) UW9 ( d31, d144 );
  not	#(1.000) UW10 ( d24, d140 );
  not	#(1.000) UW11 ( d17, d136 );
  not	#(1.000) UW12 ( d10, d132 );
  not	#(1.000) UW13 ( d109, d107 );
  not	#(1.000) UW14 ( d98, d96 );
  not	#(1.000) UW15 ( d87, d85 );
  not	#(1.000) UW16 ( d73, d71 );
  not	#(1.000) UW17 ( d120, d118 );
  nor	#(1.000) UW18 ( f2, d50, d51 );
  and	#(1.000) UW19 ( d51, d52, d53 );
  nor	#(1.000) UW20 ( d50, d52, d53 );
  nand	#(1.000) UW21 ( d53, d54, d55 );
  nor	#(1.000) UW22 ( f3, d43, d44 );
  and	#(1.000) UW23 ( d44, d45, d46 );
  nor	#(1.000) UW24 ( d43, d45, d46 );
  nand	#(1.000) UW25 ( d46, d47, d48 );
  nor	#(1.000) UW26 ( f4, d36, d37 );
  and	#(1.000) UW27 ( d37, d38, d39 );
  nor	#(1.000) UW28 ( d36, d38, d39 );
  nand	#(1.000) UW29 ( d39, d40, d41 );
  nor	#(1.000) UW30 ( f5, d29, d30 );
  and	#(1.000) UW31 ( d30, d31, d32 );
  nor	#(1.000) UW32 ( d29, d31, d32 );
  nand	#(1.000) UW33 ( d32, d33, d34 );
  nor	#(1.000) UW34 ( f6, d22, d23 );
  and	#(1.000) UW35 ( d23, d24, d25 );
  nor	#(1.000) UW36 ( d22, d24, d25 );
  nand	#(1.000) UW37 ( d25, d26, d27 );
  nor	#(1.000) UW38 ( f7, d15, d16 );
  and	#(1.000) UW39 ( d16, d17, d18 );
  nor	#(1.000) UW40 ( d15, d17, d18 );
  nand	#(1.000) UW41 ( d18, d19, d20 );
  nor	#(1.000) UW42 ( f8, d8, d9 );
  and	#(1.000) UW43 ( d9, d10, d11 );
  nor	#(1.000) UW44 ( d8, d10, d11 );
  nand	#(1.000) UW45 ( d11, d12, d13 );
  nor	#(1.000) UW46 ( f9, d1, d2 );
  and	#(1.000) UW47 ( d2, d3, d4 );
  nor	#(1.000) UW48 ( d1, d3, d4 );
  nand	#(1.000) UW49 ( d4, d5, d6 );
  nor	#(1.000) UW50 ( f10, d121, d122 );
  and	#(1.000) UW51 ( d122, d120, d123 );
  nor	#(1.000) UW52 ( d121, d120, d123 );
  nand	#(1.000) UW53 ( d123, d124, d125 );
  nor	#(1.000) UW54 ( f11, d110, d111 );
  and	#(1.000) UW55 ( d111, d109, d112 );
  nor	#(1.000) UW56 ( d110, d109, d112 );
  nand	#(1.000) UW57 ( d112, d113, d114 );
  nor	#(1.000) UW58 ( f12, d99, d100 );
  and	#(1.000) UW59 ( d100, d98, d101 );
  nor	#(1.000) UW60 ( d99, d98, d101 );
  nand	#(1.000) UW61 ( d101, d102, d103 );
  nor	#(1.000) UW62 ( f13, d88, d89 );
  and	#(1.000) UW63 ( d89, d87, d90 );
  nor	#(1.000) UW64 ( d88, d87, d90 );
  nand	#(1.000) UW65 ( d90, d91, d92 );
  nor	#(1.000) UW66 ( f14, d77, d78 );
  and	#(1.000) UW67 ( d78, d73, d79 );
  nor	#(1.000) UW68 ( d77, d73, d79 );
  nand	#(1.000) UW69 ( d79, d80, d81 );
  nor	#(1.000) UW70 ( f15, d64, d65 );
  and	#(1.000) UW71 ( d65, d66, d67 );
  nor	#(1.000) UW72 ( d64, d67, d66 );
  nand	#(1.000) UW73 ( d66, d68, d69 );
  nand	#(1.000) UW74 ( f1, d57, d58 );
  or	#(1.000) UW75 ( d58, d59, d60 );
  nand	#(1.000) UW76 ( d57, d59, d60 );
  nand	#(1.000) UW77 ( d59, d61, d62 );
  nand	#(1.000) UW78 ( d3, d129, d130 );
  nand	#(1.000) UW79 ( d129, c8, d10 );
  nand	#(1.000) UW80 ( d130, e8, d131 );
  nand	#(1.000) UW81 ( d131, d132, d14 );
  and	#(1.000) UW82 ( d156, d157, d158 );
  nand	#(1.000) UW83 ( d158, e1, d159 );
  nand	#(1.000) UW84 ( d157, c1, d160 );
  nand	#(1.000) UW85 ( d159, d63, d60 );
  and	#(1.000) UW86 ( d152, d153, d154 );
  nand	#(1.000) UW87 ( d153, c2, d52 );
  nand	#(1.000) UW88 ( d154, e2, d155 );
  nand	#(1.000) UW89 ( d155, d156, d56 );
  and	#(1.000) UW90 ( d148, d149, d150 );
  nand	#(1.000) UW91 ( d149, c3, d45 );
  nand	#(1.000) UW92 ( d150, e3, d151 );
  nand	#(1.000) UW93 ( d151, d152, d49 );
  and	#(1.000) UW94 ( d144, d145, d146 );
  nand	#(1.000) UW95 ( d145, c4, d38 );
  nand	#(1.000) UW96 ( d146, e4, d147 );
  nand	#(1.000) UW97 ( d147, d148, d42 );
  and	#(1.000) UW98 ( d107, d115, d116 );
  nand	#(1.000) UW99 ( d115, c10, d120 );
  nand	#(1.000) UW100 ( d116, e10, d117 );
  nand	#(1.000) UW101 ( d117, d118, d119 );
  and	#(1.000) UW102 ( d140, d141, d142 );
  nand	#(1.000) UW103 ( d141, c5, d31 );
  nand	#(1.000) UW104 ( d142, e5, d143 );
  nand	#(1.000) UW105 ( d143, d144, d35 );
  and	#(1.000) UW106 ( d96, d104, d105 );
  nand	#(1.000) UW107 ( d104, c11, d109 );
  nand	#(1.000) UW108 ( d105, e11, d106 );
  nand	#(1.000) UW109 ( d106, d107, d108 );
  and	#(1.000) UW110 ( d136, d137, d138 );
  nand	#(1.000) UW111 ( d137, c6, d24 );
  nand	#(1.000) UW112 ( d138, e6, d139 );
  nand	#(1.000) UW113 ( d139, d140, d28 );
  and	#(1.000) UW114 ( d85, d93, d94 );
  nand	#(1.000) UW115 ( d93, c12, d98 );
  nand	#(1.000) UW116 ( d94, e12, d95 );
  nand	#(1.000) UW117 ( d95, d96, d97 );
  and	#(1.000) UW118 ( d132, d133, d134 );
  nand	#(1.000) UW119 ( d133, c7, d17 );
  nand	#(1.000) UW120 ( d134, e7, d135 );
  nand	#(1.000) UW121 ( d135, d136, d21 );
  and	#(1.000) UW122 ( d71, d82, d83 );
  nand	#(1.000) UW123 ( d82, c13, d87 );
  nand	#(1.000) UW124 ( d83, e13, d84 );
  nand	#(1.000) UW125 ( d84, d85, d86 );
  and	#(1.000) UW126 ( d118, d126, d127 );
  nand	#(1.000) UW127 ( d127, e9, d128 );
  nand	#(1.000) UW128 ( d126, c9, d3 );
  or	#(1.000) UW129 ( d128, d3, c9 );
  nand	#(1.000) UW130 ( d67, d74, d75 );
  or	#(1.000) UW131 ( d74, d76, e15 );
  nand	#(1.000) UW132 ( d75, e15, d76 );
  not	#(1.000) UW133 ( d76, c15 );
  nand	#(1.000) UW134 ( d55, e2, d56 );
  nand	#(1.000) UW135 ( d48, e3, d49 );
  nand	#(1.000) UW136 ( d41, e4, d42 );
  nand	#(1.000) UW137 ( d34, e5, d35 );
  nand	#(1.000) UW138 ( d27, e6, d28 );
  nand	#(1.000) UW139 ( d20, e7, d21 );
  nand	#(1.000) UW140 ( d13, e8, d14 );
  nand	#(1.000) UW141 ( d125, e10, d119 );
  nand	#(1.000) UW142 ( d114, e11, d108 );
  nand	#(1.000) UW143 ( d103, e12, d97 );
  nand	#(1.000) UW144 ( d92, e13, d86 );
  nand	#(1.000) UW145 ( d81, e14, d72 );
  nand	#(1.000) UW146 ( d62, e1, d63 );
  nand	#(1.000) UW147 ( d69, e14, d70 );
  nand	#(1.000) UW148 ( d70, d71, d72 );
  nand	#(1.000) UW149 ( d68, c14, d73 );
  not	#(1.000) UW150 ( d56, c2 );
  not	#(1.000) UW151 ( d49, c3 );
  not	#(1.000) UW152 ( d42, c4 );
  not	#(1.000) UW153 ( d35, c5 );
  not	#(1.000) UW154 ( d28, c6 );
  not	#(1.000) UW155 ( d21, c7 );
  not	#(1.000) UW156 ( d14, c8 );
  not	#(1.000) UW157 ( d119, c10 );
  not	#(1.000) UW158 ( d108, c11 );
  not	#(1.000) UW159 ( d97, c12 );
  not	#(1.000) UW160 ( d86, c13 );
  not	#(1.000) UW161 ( d72, c14 );
  nand	#(1.000) UW162 ( d6, e9, d7 );
  not	#(1.000) UW163 ( d63, c1 );
  not	#(1.000) UW164 ( d161, e0 );
  not	#(1.000) UW165 ( d162, c0 );
  nand	#(1.000) UW166 ( f0, d163, d164 );
  nand	#(1.000) UW167 ( d163, c0, d161 );
  nand	#(1.000) UW168 ( d164, e0, d162 );
  or	#(1.000) UW169 ( d61, d63, e1 );
  or	#(1.000) UW170 ( d54, d56, e2 );
  or	#(1.000) UW171 ( d47, d49, e3 );
  or	#(1.000) UW172 ( d40, d42, e4 );
  or	#(1.000) UW173 ( d33, d35, e5 );
  or	#(1.000) UW174 ( d26, d28, e6 );
  or	#(1.000) UW175 ( d19, d21, e7 );
  or	#(1.000) UW176 ( d12, d14, e8 );
  or	#(1.000) UW177 ( d5, d7, e9 );
  or	#(1.000) UW178 ( d124, d119, e10 );
  or	#(1.000) UW179 ( d113, d108, e11 );
  or	#(1.000) UW180 ( d102, d97, e12 );
  or	#(1.000) UW181 ( d91, d86, e13 );
  or	#(1.000) UW182 ( d80, d72, e14 );
  not	#(1.000) UW183 ( d7, c9 );
  
  

   endmodule
  
  

          
          
          
          
          
          
          
          
          
         